`timescale 1ns / 1ps

module DataPath_tb;

    reg clk;
    reg reset;
    wire [3:0] out;
    DataPath uut (
        .clk(clk),
        .reset(reset),
        .out_1(out)
    );

    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    initial begin
    reset = 1;

    #10;
    reset = 0;
    #200;
        $finish;
end

endmodule